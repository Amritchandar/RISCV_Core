module control_store(
    input [10:0] address,
    output [16:0] control_signals
);


reg [16:0] rom[0:2062];
assign control_signals = rom[address];
initial begin
    rom[11'b01101110000] = 17'b11010100000000001;
    rom[11'b01101110001] = 17'b11010100000000001;
    rom[11'b01101110010] = 17'b11010100000000001;
    rom[11'b01101110011] = 17'b11010100000000001;
    rom[11'b01101110100] = 17'b11010100000000001;
    rom[11'b01101110101] = 17'b11010100000000001;
    rom[11'b01101110110] = 17'b11010100000000001;
    rom[11'b01101110111] = 17'b11010100000000001;
    rom[11'b01101111000] = 17'b11010100000000001;
    rom[11'b01101111001] = 17'b11010100000000001;
    rom[11'b01101111010] = 17'b11010100000000001;
    rom[11'b01101111011] = 17'b11010100000000001;
    rom[11'b01101111100] = 17'b11010100000000001;
    rom[11'b01101111101] = 17'b11010100000000001;
    rom[11'b01101111110] = 17'b11010100000000001;
    rom[11'b01101111111] = 17'b11010100000000001;
    rom[11'b00101110000] = 17'b11010110000000001;
    rom[11'b00101110001] = 17'b11010110000000001;
    rom[11'b00101110010] = 17'b11010110000000001;
    rom[11'b00101110011] = 17'b11010110000000001;
    rom[11'b00101110100] = 17'b11010110000000001;
    rom[11'b00101110101] = 17'b11010110000000001;
    rom[11'b00101110110] = 17'b11010110000000001;
    rom[11'b00101110111] = 17'b11010110000000001;
    rom[11'b00101111000] = 17'b11010110000000001;
    rom[11'b00101111001] = 17'b11010110000000001;
    rom[11'b00101111010] = 17'b11010110000000001;
    rom[11'b00101111011] = 17'b11010110000000001;
    rom[11'b00101111100] = 17'b11010110000000001;
    rom[11'b00101111101] = 17'b11010110000000001;
    rom[11'b00101111110] = 17'b11010110000000001;
    rom[11'b00101111111] = 17'b11010110000000001;
    rom[11'b11011110000] = 17'b11011000000000001;
    rom[11'b11011110001] = 17'b11011000000000001;
    rom[11'b11011110010] = 17'b11011000000000001;
    rom[11'b11011110011] = 17'b11011000000000001;
    rom[11'b11011110100] = 17'b11011000000000001;
    rom[11'b11011110101] = 17'b11011000000000001;
    rom[11'b11011110110] = 17'b11011000000000001;
    rom[11'b11011110111] = 17'b11011000000000001;
    rom[11'b11011111000] = 17'b11011000000000001;
    rom[11'b11011111001] = 17'b11011000000000001;
    rom[11'b11011111010] = 17'b11011000000000001;
    rom[11'b11011111011] = 17'b11011000000000001;
    rom[11'b11011111100] = 17'b11011000000000001;
    rom[11'b11011111101] = 17'b11011000000000001;
    rom[11'b11011111110] = 17'b11011000000000001;
    rom[11'b11011111111] = 17'b11011000000000001;
    rom[11'b11001110000] = 17'b11011000000000001;
    rom[11'b11001110001] = 17'b11011000000000001;
    rom[11'b11000110000] = 17'b00011010000000000;
    rom[11'b11000110001] = 17'b00011010000000000;
    rom[11'b11000110010] = 17'b00111010000000000;
    rom[11'b11000110011] = 17'b00111010000000000;
    rom[11'b11000111000] = 17'b01011010000000000;
    rom[11'b11000111001] = 17'b01011010000000000;
    rom[11'b11000111010] = 17'b01111010000000000;
    rom[11'b11000111011] = 17'b01111010000000000;
    rom[11'b11000111100] = 17'b10011010000000000;
    rom[11'b11000111101] = 17'b10011010000000000;
    rom[11'b11000111110] = 17'b10111010000000000;
    rom[11'b11000111111] = 17'b10111010000000000;
    rom[11'b00000110000] = 17'b11011010000000011;
    rom[11'b00000110001] = 17'b11011010000000011;
    rom[11'b00000110010] = 17'b11011010000000111;
    rom[11'b00000110011] = 17'b11011010000000111;
    rom[11'b00000110100] = 17'b11011010000001011;
    rom[11'b00000110101] = 17'b11011010000001011;
    rom[11'b00000111000] = 17'b11011010000001111;
    rom[11'b00000111001] = 17'b11011010000001111;
    rom[11'b00000111010] = 17'b11011010000010011;
    rom[11'b00000111011] = 17'b11011010000010011;
    rom[11'b01000110000] = 17'b11010100000100000;
    rom[11'b01000110001] = 17'b11010100000100000;
    rom[11'b01000110010] = 17'b11010100000100000;
    rom[11'b01000110011] = 17'b11010100000100000;
    rom[11'b01000110100] = 17'b11010100000100000;
    rom[11'b01000110101] = 17'b11010100000100000;
    rom[11'b00100110000] = 17'b11000000000000001;
    rom[11'b00100110001] = 17'b11000000000000001;
    rom[11'b00100110100] = 17'b11000110000000001;
    rom[11'b00100110101] = 17'b11000110000000001;
    rom[11'b00100110110] = 17'b11001000000000001;
    rom[11'b00100110111] = 17'b11001000000000001;
    rom[11'b00100111000] = 17'b11001010000000001;
    rom[11'b00100111001] = 17'b11001010000000001;
    rom[11'b00100111100] = 17'b11010000000000001;
    rom[11'b00100111101] = 17'b11010000000000001;
    rom[11'b00100111110] = 17'b11010010000000001;
    rom[11'b00100111111] = 17'b11010010000000001;
    rom[11'b00100110010] = 17'b11000100000000001;
    rom[11'b00100111010] = 17'b11001100000000001;
    rom[11'b00100111011] = 17'b11001110000000001;
    rom[11'b01100110000] = 17'b11000000000000001;
    rom[11'b01100110001] = 17'b11000010000000001;
    rom[11'b01100110010] = 17'b11000100000000001;
    rom[11'b01100110100] = 17'b11000110000000001;
    rom[11'b01100110110] = 17'b11001000000000001;
    rom[11'b01100111000] = 17'b11001010000000001;
    rom[11'b01100111010] = 17'b11001100000000001;
    rom[11'b01100111011] = 17'b11001110000000001;
    rom[11'b01100111100] = 17'b11010000000000001;
    rom[11'b01100111110] = 17'b11010010000000001;
    rom[11'b00000111100] = 17'b11011010000010111;
    rom[11'b00000111101] = 17'b11011010000010111;
    rom[11'b00000110110] = 17'b11011010000011011;
    rom[11'b01000110110] = 17'b11010100000100000;
    rom[11'b01000110111] = 17'b11010100000100000;
    rom[11'b00110110000] = 17'b11000000000000001;
    rom[11'b00110110001] = 17'b11000000000000001;
    rom[11'b00110110010] = 17'b11000100000000001;
    rom[11'b00110111010] = 17'b11001100000000001;
    rom[11'b00110111011] = 17'b11001110000000001;
    rom[11'b01110110000] = 17'b11000000000000001;
    rom[11'b01110110001] = 17'b11000010000000001;
    rom[11'b01110110010] = 17'b11000100000000001;
    rom[11'b01110111010] = 17'b11001100000000001;
    rom[11'b01110111011] = 17'b11001110000000001;
    rom[11'b01100110000] = 17'b11011011000000001;
    rom[11'b01100110010] = 17'b11011011001000001;
    rom[11'b01100110100] = 17'b11011011010000001;
    rom[11'b01100110110] = 17'b11011011011000001;
    rom[11'b01100111000] = 17'b11011011100000001;
    rom[11'b01100111010] = 17'b11011011101000001;
    rom[11'b01100111100] = 17'b11011011110000001;
    rom[11'b01100111110] = 17'b11011011101000001;
    rom[11'b01110110000] = 17'b11011011000000001;
    rom[11'b01110111000] = 17'b11011011100000001;
    rom[11'b01110111010] = 17'b11011011101000001;
    rom[11'b01110111100] = 17'b11011011110000001;
    rom[11'b01110111110] = 17'b11011011111000001;
end
endmodule