module control_store(
    input [11:0] address,
    output [18:0] control_signals
);

reg [18:0] rom[0:8000];

assign control_signals = rom[address];
initial begin
    // LUI
    rom[12'b011011100000] = 19'b0011110100000000001;
    rom[12'b011011100001] = 19'b0011110100000000001;
    rom[12'b011011100010] = 19'b0011110100000000001;
    rom[12'b011011100011] = 19'b0011110100000000001;
    rom[12'b011011100100] = 19'b0011110100000000001;
    rom[12'b011011100101] = 19'b0011110100000000001;
    rom[12'b011011100110] = 19'b0011110100000000001;
    rom[12'b011011100111] = 19'b0011110100000000001;
    rom[12'b011011101000] = 19'b0011110100000000001;
    rom[12'b011011101001] = 19'b0011110100000000001;
    rom[12'b011011101010] = 19'b0011110100000000001;
    rom[12'b011011101011] = 19'b0011110100000000001;
    rom[12'b011011101100] = 19'b0011110100000000001;
    rom[12'b011011101101] = 19'b0011110100000000001;
    rom[12'b011011101110] = 19'b0011110100000000001;
    rom[12'b011011101111] = 19'b0011110100000000001;
    rom[12'b011011110000] = 19'b0011110100000000001;
    rom[12'b011011110001] = 19'b0011110100000000001;
    rom[12'b011011110010] = 19'b0011110100000000001;
    rom[12'b011011110011] = 19'b0011110100000000001;
    rom[12'b011011110100] = 19'b0011110100000000001;
    rom[12'b011011110101] = 19'b0011110100000000001;
    rom[12'b011011110110] = 19'b0011110100000000001;
    rom[12'b011011110111] = 19'b0011110100000000001;
    rom[12'b011011111000] = 19'b0011110100000000001;
    rom[12'b011011111001] = 19'b0011110100000000001;
    rom[12'b011011111010] = 19'b0011110100000000001;
    rom[12'b011011111011] = 19'b0011110100000000001;
    rom[12'b011011111100] = 19'b0011110100000000001;
    rom[12'b011011111101] = 19'b0011110100000000001;
    rom[12'b011011111110] = 19'b0011110100000000001;
    rom[12'b011011111111] = 19'b0011110100000000001;
    // AUIPC
    rom[12'b001011100000] = 19'b0011110110000000001;
    rom[12'b001011100001] = 19'b0011110110000000001;
    rom[12'b001011100010] = 19'b0011110110000000001;
    rom[12'b001011100011] = 19'b0011110110000000001;
    rom[12'b001011100100] = 19'b0011110110000000001;
    rom[12'b001011100101] = 19'b0011110110000000001;
    rom[12'b001011100110] = 19'b0011110110000000001;
    rom[12'b001011100111] = 19'b0011110110000000001;
    rom[12'b001011101000] = 19'b0011110110000000001;
    rom[12'b001011101001] = 19'b0011110110000000001;
    rom[12'b001011101010] = 19'b0011110110000000001;
    rom[12'b001011101011] = 19'b0011110110000000001;
    rom[12'b001011101100] = 19'b0011110110000000001;
    rom[12'b001011101101] = 19'b0011110110000000001;
    rom[12'b001011101110] = 19'b0011110110000000001;
    rom[12'b001011101111] = 19'b0011110110000000001;
    rom[12'b001011110000] = 19'b0011110110000000001;
    rom[12'b001011110001] = 19'b0011110110000000001;
    rom[12'b001011110010] = 19'b0011110110000000001;
    rom[12'b001011110011] = 19'b0011110110000000001;
    rom[12'b001011110100] = 19'b0011110110000000001;
    rom[12'b001011110101] = 19'b0011110110000000001;
    rom[12'b001011110110] = 19'b0011110110000000001;
    rom[12'b001011110111] = 19'b0011110110000000001;
    rom[12'b001011111000] = 19'b0011110110000000001;
    rom[12'b001011111001] = 19'b0011110110000000001;
    rom[12'b001011111010] = 19'b0011110110000000001;
    rom[12'b001011111011] = 19'b0011110110000000001;
    rom[12'b001011111100] = 19'b0011110110000000001;
    rom[12'b001011111101] = 19'b0011110110000000001;
    rom[12'b001011111110] = 19'b0011110110000000001;
    rom[12'b001011111111] = 19'b0011110110000000001;
    // JAL
    rom[12'b110111100000] = 19'b0011011000000000001;
    rom[12'b110111100001] = 19'b0011011000000000001;
    rom[12'b110111100010] = 19'b0011011000000000001;
    rom[12'b110111100011] = 19'b0011011000000000001;
    rom[12'b110111100100] = 19'b0011011000000000001;
    rom[12'b110111100101] = 19'b0011011000000000001;
    rom[12'b110111100110] = 19'b0011011000000000001;
    rom[12'b110111100111] = 19'b0011011000000000001;
    rom[12'b110111101000] = 19'b0011011000000000001;
    rom[12'b110111101001] = 19'b0011011000000000001;
    rom[12'b110111101010] = 19'b0011011000000000001;
    rom[12'b110111101011] = 19'b0011011000000000001;
    rom[12'b110111101100] = 19'b0011011000000000001;
    rom[12'b110111101101] = 19'b0011011000000000001;
    rom[12'b110111101110] = 19'b0011011000000000001;
    rom[12'b110111101111] = 19'b0011011000000000001;
    rom[12'b110111110000] = 19'b0011011000000000001;
    rom[12'b110111110001] = 19'b0011011000000000001;
    rom[12'b110111110010] = 19'b0011011000000000001;
    rom[12'b110111110011] = 19'b0011011000000000001;
    rom[12'b110111110100] = 19'b0011011000000000001;
    rom[12'b110111110101] = 19'b0011011000000000001;
    rom[12'b110111110110] = 19'b0011011000000000001;
    rom[12'b110111110111] = 19'b0011011000000000001;
    rom[12'b110111111000] = 19'b0011011000000000001;
    rom[12'b110111111001] = 19'b0011011000000000001;
    rom[12'b110111111010] = 19'b0011011000000000001;
    rom[12'b110111111011] = 19'b0011011000000000001;
    rom[12'b110111111100] = 19'b0011011000000000001;
    rom[12'b110111111101] = 19'b0011011000000000001;
    rom[12'b110111111110] = 19'b0011011000000000001;
    rom[12'b110111111111] = 19'b0011011000000000001;
    // JALR
    rom[12'b110011100000] = 19'b0011011000000000001;
    rom[12'b110011100001] = 19'b0011011000000000001;
    rom[12'b110011100010] = 19'b0011011000000000001;
    rom[12'b110011100011] = 19'b0011011000000000001;
    // BEQ
    rom[12'b110001100000] = 19'b0000011010000000000;
    rom[12'b110001100001] = 19'b0000011010000000000;
    rom[12'b110001100010] = 19'b0000011010000000000;
    rom[12'b110001100011] = 19'b0000011010000000000;
    // BNE
    rom[12'b110001100100] = 19'b0000111010000000000;
    rom[12'b110001100101] = 19'b0000111010000000000;
    rom[12'b110001100110] = 19'b0000111010000000000;
    rom[12'b110001100111] = 19'b0000111010000000000;
    // BLT
    rom[12'b110001110000] = 19'b0001011010000000000;
    rom[12'b110001110001] = 19'b0001011010000000000;
    rom[12'b110001110010] = 19'b0001011010000000000;
    rom[12'b110001110011] = 19'b0001011010000000000;
    // BGE
    rom[12'b110001110100] = 19'b0001111010000000000;
    rom[12'b110001110101] = 19'b0001111010000000000;
    rom[12'b110001110110] = 19'b0001111010000000000;
    rom[12'b110001110111] = 19'b0001111010000000000;
    // BLTU
    rom[12'b110001111000] = 19'b0010011010000000000;
    rom[12'b110001111001] = 19'b0010011010000000000;
    rom[12'b110001111010] = 19'b0010011010000000000;
    rom[12'b110001111011] = 19'b0010011010000000000;
    // BGEU
    rom[12'b110001111100] = 19'b0010111010000000000;
    rom[12'b110001111101] = 19'b0010111010000000000;
    rom[12'b110001111110] = 19'b0010111010000000000;
    rom[12'b110001111111] = 19'b0010111010000000000;
    // LB
    rom[12'b000001100000] = 19'b0011111010000000011;
    rom[12'b000001100001] = 19'b0011111010000000011;
    rom[12'b000001100010] = 19'b0011111010000000011;
    rom[12'b000001100011] = 19'b0011111010000000011;
    // LH
    rom[12'b000001100100] = 19'b0011111010000000111;
    rom[12'b000001100101] = 19'b0011111010000000111;
    rom[12'b000001100110] = 19'b0011111010000000111;
    rom[12'b000001100111] = 19'b0011111010000000111;
    // LW
    rom[12'b000001101000] = 19'b0011111010000001011;
    rom[12'b000001101001] = 19'b0011111010000001011;
    rom[12'b000001101010] = 19'b0011111010000001011;
    rom[12'b000001101011] = 19'b0011111010000001011;
    // LBU
    rom[12'b000001110000] = 19'b0011111010000001111;
    rom[12'b000001110001] = 19'b0011111010000001111;
    rom[12'b000001110010] = 19'b0011111010000001111;
    rom[12'b000001110011] = 19'b0011111010000001111;
    // LHU
    rom[12'b000001110100] = 19'b0011111010000010011;
    rom[12'b000001110101] = 19'b0011111010000010011;
    rom[12'b000001110110] = 19'b0011111010000010011;
    rom[12'b000001110111] = 19'b0011111010000010011;
    // SB
    rom[12'b010001100000] = 19'b0011110100000100000;
    rom[12'b010001100001] = 19'b0011110100000100000;
    rom[12'b010001100010] = 19'b0011110100000100000;
    rom[12'b010001100011] = 19'b0011110100000100000;
    // SH
    rom[12'b010001100100] = 19'b0011110100000100000;
    rom[12'b010001100101] = 19'b0011110100000100000;
    rom[12'b010001100110] = 19'b0011110100000100000;
    rom[12'b010001100111] = 19'b0011110100000100000;
    // SW
    rom[12'b010001101000] = 19'b0011110100000100000;
    rom[12'b010001101001] = 19'b0011110100000100000;
    rom[12'b010001101010] = 19'b0011110100000100000;
    rom[12'b010001101011] = 19'b0011110100000100000;
    // ADDI
    rom[12'b001001100000] = 19'b0011100000000000001;
    rom[12'b001001100001] = 19'b0011100000000000001;
    rom[12'b001001100010] = 19'b0011100000000000001;
    rom[12'b001001100011] = 19'b0011100000000000001;
    // SLTI
    rom[12'b001001101000] = 19'b0011100110000000001;
    rom[12'b001001101001] = 19'b0011100110000000001;
    rom[12'b001001101010] = 19'b0011100110000000001;
    rom[12'b001001101011] = 19'b0011100110000000001;
    // SLTIU
    rom[12'b001001101100] = 19'b0011101000000000001;
    rom[12'b001001101101] = 19'b0011101000000000001;
    rom[12'b001001101110] = 19'b0011101000000000001;
    rom[12'b001001101111] = 19'b0011101000000000001;
    // XORI
    rom[12'b001001110000] = 19'b0011101010000000001;
    rom[12'b001001110001] = 19'b0011101010000000001;
    rom[12'b001001110010] = 19'b0011101010000000001;
    rom[12'b001001110011] = 19'b0011101010000000001;
    // ORI
    rom[12'b001001111000] = 19'b0011110000000000001;
    rom[12'b001001111001] = 19'b0011110000000000001;
    rom[12'b001001111010] = 19'b0011110000000000001;
    rom[12'b001001111011] = 19'b0011110000000000001;
    // ANDI
    rom[12'b001001111100] = 19'b0011110010000000001;
    rom[12'b001001111101] = 19'b0011110010000000001;
    rom[12'b001001111110] = 19'b0011110010000000001;
    rom[12'b001001111111] = 19'b0011110010000000001;
    // SLLI
    rom[12'b001001100100] = 19'b0011100100000000001;
    // SRLI
    rom[12'b001001110100] = 19'b0011101100000000001;
    // SRAI
    rom[12'b001001110110] = 19'b0011101110000000001;
    // ADD
    rom[12'b011001100000] = 19'b0011100000000000001;
    // SUB
    rom[12'b011001100010] = 19'b0011100010000000001;
    // SLL
    rom[12'b011001100100] = 19'b0011100100000000001;
    // SLT
    rom[12'b011001101000] = 19'b0011100110000000001;
    // SLTU
    rom[12'b011001101100] = 19'b0011101000000000001;
    // XOR
    rom[12'b011001110000] = 19'b0011101010000000001;
    // SRL
    rom[12'b011001110100] = 19'b0011101100000000001;
    // SRA
    rom[12'b011001110110] = 19'b0011101110000000001;
    // OR
    rom[12'b011001111000] = 19'b0011110000000000001;
    // AND
    rom[12'b011001111100] = 19'b0011110010000000001;
    // LWU
    rom[12'b000001111000] = 19'b0011111010000010111;
    rom[12'b000001111001] = 19'b0011111010000010111;
    rom[12'b000001111010] = 19'b0011111010000010111;
    rom[12'b000001111011] = 19'b0011111010000010111;
    // LD
    rom[12'b000001101100] = 19'b0011111010000011011;
    rom[12'b000001101101] = 19'b0011111010000011011;
    rom[12'b000001101110] = 19'b0011111010000011011;
    rom[12'b000001101111] = 19'b0011111010000011011;
    // SD
    rom[12'b010001101100] = 19'b0011110100000100000;
    rom[12'b010001101101] = 19'b0011110100000100000;
    rom[12'b010001101110] = 19'b0011110100000100000;
    rom[12'b010001101111] = 19'b0011110100000100000;
    // ADDIW
    rom[12'b001101100000] = 19'b0111100000000000001;
    rom[12'b001101100001] = 19'b0111100000000000001;
    rom[12'b001101100010] = 19'b0111100000000000001;
    rom[12'b001101100011] = 19'b0111100000000000001;
    // SLLIW
    rom[12'b001101100100] = 19'b0111100100000000001;
    // SRLIW
    rom[12'b001101110100] = 19'b0111101100000000001;
    // SRAIW
    rom[12'b001101110110] = 19'b0111101110000000001;
    // ADDW
    rom[12'b011101100000] = 19'b0111100000000000001;
    // SUBW
    rom[12'b011101100010] = 19'b0111100010000000001;
    // SLLW
    rom[12'b011101100100] = 19'b0111100100000000001;
    // SRLW
    rom[12'b011101110100] = 19'b0111101100000000001;
    // SRAW
    rom[12'b011101110110] = 19'b0111101110000000001;
    // MUL
    rom[12'b011001100001] = 19'b0011111011000000001;
    // MULH
    rom[12'b011001100101] = 19'b0011111011001000001;
    // MULHSU
    rom[12'b011001101001] = 19'b0011111011010000001;
    // MULHU
    rom[12'b011001101101] = 19'b0011111011011000001;
    // DIV
    rom[12'b011001110001] = 19'b0011111011100000001;
    // DIVU
    rom[12'b011001110101] = 19'b0011111011101000001;
    // REM
    rom[12'b011001111001] = 19'b0011111011110000001;
    // REMU
    rom[12'b011001111101] = 19'b0011111011101000001;
    // MULW
    rom[12'b011101100001] = 19'b0111111011000000001;
    // DIVW
    rom[12'b011101110001] = 19'b0111111011100000001;
    // DIVUW
    rom[12'b011101110101] = 19'b1111111011101000001;
    // REMW
    rom[12'b011101111001] = 19'b0111111011110000001;
    // REMUW
    rom[12'b011101111101] = 19'b1111111011111000001;
end
endmodule
